module bru #(
    parameter Width = 32
) (
    ports
);

endmodule
