localparam Width = 32;
