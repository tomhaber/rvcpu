package rvcpu;

typedef enum {auipc_imm, alu_imm, uimm, load_offset, store_offset, jal_offset, jalr_offset, br_offset, none} imm_type_t;

endpackage : rvcpu
