
`timescale 1ns / 1ps

module top
  (input logic clk,
   input logic reset);

sext_tb sext_tb();

endmodule
